`ifndef __OUT_TRANS__
`define __OUT_TRANS__

class out_trans extends router_trans_base;

   logic data [];

endclass

`endif
