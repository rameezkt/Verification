

// here you have to instantiate in_agent[num_port] and out_agent[num_port],router_scoreboard
// and make the required connection for the scoreboard
